//=============================================================================
// Project       : UART VIP
//=============================================================================
// Filename      : seq_pkg.sv
// Author        : Huy Nguyen
// Company       : NO
// Date          : 20-Dec-2021
//=============================================================================
// Description   : 
//
//
//
//=============================================================================
`ifndef GUARD_UART_SEQ_PKG__SV
`define GUARD_UART_SEQ_PKG__SV

package seq_pkg;
  import uvm_pkg::*;
  import uart_pkg::*;
	import ahb_pkg::*;
  // Include your file
	`include "uart_sequence.sv" 
	`include "uart_sequence_cont.sv" 
	`include "uart_sequence_cont_17.sv"
	`include "access_rsvd_sequence.sv" 

endpackage: seq_pkg

`endif


