package test_pkg;
  import uvm_pkg::*;
  import ahb_pkg::*;
  import env_pkg::*;
  import seq_pkg::*;
  import uart_regmodel_pkg::*;
	
	import uart_pkg::*;

  `include "uart_base_test.sv"

	/*--------------------------REGISTER TEST--------------------------*/
  `include "uart_reg_scan_test.sv"	
  `include "parity_error_w1c.sv"
		

	/*--------------------------OVERSAMPLING--------------------------*/
	//16x - baudrate
   `include "x16_2400.sv"
   `include "x16_4800.sv"
   `include "x16_9600.sv"
   `include "x16_19200.sv"
   `include "x16_38400.sv"
   `include "x16_76800.sv"
   `include "x16_115200.sv"
   `include "x16_230400.sv"	

	//13x - baudrate
   `include "x13_2400.sv"
   `include "x13_4800.sv"
   `include "x13_9600.sv"
   `include "x13_19200.sv"
   `include "x13_38400.sv"
   `include "x13_76800.sv"
   `include "x13_115200.sv"
   `include "x13_230400.sv"


	 /*---------------------TRANSMITTER TEST-----------------------*/
	
   `include "tx_2400_5_no_1.sv"
   `include "tx_2400_6_no_1.sv"
   `include "tx_2400_7_no_1.sv"
   `include "tx_2400_8_no_1.sv"
   `include "tx_2400_5_even_1.sv"
   `include "tx_2400_6_even_1.sv"
   `include "tx_2400_7_even_1.sv"
   `include "tx_2400_8_even_1.sv"
   `include "tx_2400_5_odd_1.sv"
   `include "tx_2400_6_odd_1.sv"
   `include "tx_2400_7_odd_1.sv"
   `include "tx_2400_8_odd_1.sv"
   `include "tx_2400_5_no_2.sv"
   `include "tx_2400_6_no_2.sv"
   `include "tx_2400_7_no_2.sv"
   `include "tx_2400_8_no_2.sv"
   `include "tx_2400_5_even_2.sv"
   `include "tx_2400_6_even_2.sv"
   `include "tx_2400_7_even_2.sv"
   `include "tx_2400_8_even_2.sv"
   `include "tx_2400_5_odd_2.sv"
   `include "tx_2400_6_odd_2.sv"
   `include "tx_2400_7_odd_2.sv"
   `include "tx_2400_8_odd_2.sv"
   `include "tx_4800_5_no_1.sv"
   `include "tx_4800_6_no_1.sv"
   `include "tx_4800_7_no_1.sv"
   `include "tx_4800_8_no_1.sv"
   `include "tx_4800_5_even_1.sv"
   `include "tx_4800_6_even_1.sv"
   `include "tx_4800_7_even_1.sv"
   `include "tx_4800_8_even_1.sv"
   `include "tx_4800_5_odd_1.sv"
   `include "tx_4800_6_odd_1.sv"
   `include "tx_4800_7_odd_1.sv"
   `include "tx_4800_8_odd_1.sv"
   `include "tx_4800_5_no_2.sv"
   `include "tx_4800_6_no_2.sv"
   `include "tx_4800_7_no_2.sv"
   `include "tx_4800_8_no_2.sv"
   `include "tx_4800_5_even_2.sv"
   `include "tx_4800_6_even_2.sv"
   `include "tx_4800_7_even_2.sv"
   `include "tx_4800_8_even_2.sv"
   `include "tx_4800_5_odd_2.sv"
   `include "tx_4800_6_odd_2.sv"
   `include "tx_4800_7_odd_2.sv"
   `include "tx_4800_8_odd_2.sv"
   `include "tx_9600_5_no_1.sv"
   `include "tx_9600_6_no_1.sv"
   `include "tx_9600_7_no_1.sv"
   `include "tx_9600_8_no_1.sv"
   `include "tx_9600_5_even_1.sv"
   `include "tx_9600_6_even_1.sv"
   `include "tx_9600_7_even_1.sv"
   `include "tx_9600_8_even_1.sv"
   `include "tx_9600_5_odd_1.sv"
   `include "tx_9600_6_odd_1.sv"
   `include "tx_9600_7_odd_1.sv"
   `include "tx_9600_8_odd_1.sv"
   `include "tx_9600_5_no_2.sv"
   `include "tx_9600_6_no_2.sv"
   `include "tx_9600_7_no_2.sv"
   `include "tx_9600_8_no_2.sv"
   `include "tx_9600_5_even_2.sv"
   `include "tx_9600_6_even_2.sv"
   `include "tx_9600_7_even_2.sv"
   `include "tx_9600_8_even_2.sv"
   `include "tx_9600_5_odd_2.sv"
   `include "tx_9600_6_odd_2.sv"
   `include "tx_9600_7_odd_2.sv"
   `include "tx_9600_8_odd_2.sv"
   `include "tx_19200_5_no_1.sv"
   `include "tx_19200_6_no_1.sv"
   `include "tx_19200_7_no_1.sv"
   `include "tx_19200_8_no_1.sv"
   `include "tx_19200_5_even_1.sv"
   `include "tx_19200_6_even_1.sv"
   `include "tx_19200_7_even_1.sv"
   `include "tx_19200_8_even_1.sv"
   `include "tx_19200_5_odd_1.sv"
   `include "tx_19200_6_odd_1.sv"
   `include "tx_19200_7_odd_1.sv"
   `include "tx_19200_8_odd_1.sv"
   `include "tx_19200_5_no_2.sv"
   `include "tx_19200_6_no_2.sv"
   `include "tx_19200_7_no_2.sv"
   `include "tx_19200_8_no_2.sv"
   `include "tx_19200_5_even_2.sv"
   `include "tx_19200_6_even_2.sv"
   `include "tx_19200_7_even_2.sv"
   `include "tx_19200_8_even_2.sv"
   `include "tx_19200_5_odd_2.sv"
   `include "tx_19200_6_odd_2.sv"
   `include "tx_19200_7_odd_2.sv"
   `include "tx_19200_8_odd_2.sv"
   `include "tx_38400_5_no_1.sv"
   `include "tx_38400_6_no_1.sv"
   `include "tx_38400_7_no_1.sv"
   `include "tx_38400_8_no_1.sv"
   `include "tx_38400_5_even_1.sv"
   `include "tx_38400_6_even_1.sv"
   `include "tx_38400_7_even_1.sv"
   `include "tx_38400_8_even_1.sv"
   `include "tx_38400_5_odd_1.sv"
   `include "tx_38400_6_odd_1.sv"
   `include "tx_38400_7_odd_1.sv"
   `include "tx_38400_8_odd_1.sv"
   `include "tx_38400_5_no_2.sv"
   `include "tx_38400_6_no_2.sv"
   `include "tx_38400_7_no_2.sv"
   `include "tx_38400_8_no_2.sv"
   `include "tx_38400_5_even_2.sv"
   `include "tx_38400_6_even_2.sv"
   `include "tx_38400_7_even_2.sv"
   `include "tx_38400_8_even_2.sv"
   `include "tx_38400_5_odd_2.sv"
   `include "tx_38400_6_odd_2.sv"
   `include "tx_38400_7_odd_2.sv"
   `include "tx_38400_8_odd_2.sv"
   `include "tx_76800_5_no_1.sv"
   `include "tx_76800_6_no_1.sv"
   `include "tx_76800_7_no_1.sv"
   `include "tx_76800_8_no_1.sv"
   `include "tx_76800_5_even_1.sv"
   `include "tx_76800_6_even_1.sv"
   `include "tx_76800_7_even_1.sv"
   `include "tx_76800_8_even_1.sv"
   `include "tx_76800_5_odd_1.sv"
   `include "tx_76800_6_odd_1.sv"
   `include "tx_76800_7_odd_1.sv"
   `include "tx_76800_8_odd_1.sv"
   `include "tx_76800_5_no_2.sv"
   `include "tx_76800_6_no_2.sv"
   `include "tx_76800_7_no_2.sv"
   `include "tx_76800_8_no_2.sv"
   `include "tx_76800_5_even_2.sv"
   `include "tx_76800_6_even_2.sv"
   `include "tx_76800_7_even_2.sv"
   `include "tx_76800_8_even_2.sv"
   `include "tx_76800_5_odd_2.sv"
   `include "tx_76800_6_odd_2.sv"
   `include "tx_76800_7_odd_2.sv"
   `include "tx_76800_8_odd_2.sv"
   `include "tx_115200_5_no_1.sv"
   `include "tx_115200_6_no_1.sv"
   `include "tx_115200_7_no_1.sv"
   `include "tx_115200_8_no_1.sv"
   `include "tx_115200_5_even_1.sv"
   `include "tx_115200_6_even_1.sv"
   `include "tx_115200_7_even_1.sv"
   `include "tx_115200_8_even_1.sv"
   `include "tx_115200_5_odd_1.sv"
   `include "tx_115200_6_odd_1.sv"
   `include "tx_115200_7_odd_1.sv"
   `include "tx_115200_8_odd_1.sv"
   `include "tx_115200_5_no_2.sv"
   `include "tx_115200_6_no_2.sv"
   `include "tx_115200_7_no_2.sv"
   `include "tx_115200_8_no_2.sv"
   `include "tx_115200_5_even_2.sv"
   `include "tx_115200_6_even_2.sv"
   `include "tx_115200_7_even_2.sv"
   `include "tx_115200_8_even_2.sv"
   `include "tx_115200_5_odd_2.sv"
   `include "tx_115200_6_odd_2.sv"
   `include "tx_115200_7_odd_2.sv"
   `include "tx_115200_8_odd_2.sv"
   `include "tx_230400_5_no_1.sv"
   `include "tx_230400_6_no_1.sv"
   `include "tx_230400_7_no_1.sv"
   `include "tx_230400_8_no_1.sv"
   `include "tx_230400_5_even_1.sv"
   `include "tx_230400_6_even_1.sv"
   `include "tx_230400_7_even_1.sv"
   `include "tx_230400_8_even_1.sv"
   `include "tx_230400_5_odd_1.sv"
   `include "tx_230400_6_odd_1.sv"
   `include "tx_230400_7_odd_1.sv"
   `include "tx_230400_8_odd_1.sv"
   `include "tx_230400_5_no_2.sv"
   `include "tx_230400_6_no_2.sv"
   `include "tx_230400_7_no_2.sv"
   `include "tx_230400_8_no_2.sv"
   `include "tx_230400_5_even_2.sv"
   `include "tx_230400_6_even_2.sv"
   `include "tx_230400_7_even_2.sv"
   `include "tx_230400_8_even_2.sv"
   `include "tx_230400_5_odd_2.sv"
   `include "tx_230400_6_odd_2.sv"
   `include "tx_230400_7_odd_2.sv"
   `include "tx_230400_8_odd_2.sv"


	 /*---------------------RECEIVER TEST-----------------------*/
   `include "rx_2400_5_no_1.sv"
   `include "rx_2400_6_no_1.sv"
   `include "rx_2400_7_no_1.sv"
   `include "rx_2400_8_no_1.sv"
   `include "rx_2400_5_even_1.sv"
   `include "rx_2400_6_even_1.sv"
   `include "rx_2400_7_even_1.sv"
   `include "rx_2400_8_even_1.sv"
   `include "rx_2400_5_odd_1.sv"
   `include "rx_2400_6_odd_1.sv"
   `include "rx_2400_7_odd_1.sv"
   `include "rx_2400_8_odd_1.sv"
   `include "rx_2400_5_no_2.sv"
   `include "rx_2400_6_no_2.sv"
   `include "rx_2400_7_no_2.sv"
   `include "rx_2400_8_no_2.sv"
   `include "rx_2400_5_even_2.sv"
   `include "rx_2400_6_even_2.sv"
   `include "rx_2400_7_even_2.sv"
   `include "rx_2400_8_even_2.sv"
   `include "rx_2400_5_odd_2.sv"
   `include "rx_2400_6_odd_2.sv"
   `include "rx_2400_7_odd_2.sv"
   `include "rx_2400_8_odd_2.sv"
   `include "rx_4800_5_no_1.sv"
   `include "rx_4800_6_no_1.sv"
   `include "rx_4800_7_no_1.sv"
   `include "rx_4800_8_no_1.sv"
   `include "rx_4800_5_even_1.sv"
   `include "rx_4800_6_even_1.sv"
   `include "rx_4800_7_even_1.sv"
   `include "rx_4800_8_even_1.sv"
   `include "rx_4800_5_odd_1.sv"
   `include "rx_4800_6_odd_1.sv"
   `include "rx_4800_7_odd_1.sv"
   `include "rx_4800_8_odd_1.sv"
   `include "rx_4800_5_no_2.sv"
   `include "rx_4800_6_no_2.sv"
   `include "rx_4800_7_no_2.sv"
   `include "rx_4800_8_no_2.sv"
   `include "rx_4800_5_even_2.sv"
   `include "rx_4800_6_even_2.sv"
   `include "rx_4800_7_even_2.sv"
   `include "rx_4800_8_even_2.sv"
   `include "rx_4800_5_odd_2.sv"
   `include "rx_4800_6_odd_2.sv"
   `include "rx_4800_7_odd_2.sv"
   `include "rx_4800_8_odd_2.sv"
   `include "rx_9600_5_no_1.sv"
   `include "rx_9600_6_no_1.sv"
   `include "rx_9600_7_no_1.sv"
   `include "rx_9600_8_no_1.sv"
   `include "rx_9600_5_even_1.sv"
   `include "rx_9600_6_even_1.sv"
   `include "rx_9600_7_even_1.sv"
   `include "rx_9600_8_even_1.sv"
   `include "rx_9600_5_odd_1.sv"
   `include "rx_9600_6_odd_1.sv"
   `include "rx_9600_7_odd_1.sv"
   `include "rx_9600_8_odd_1.sv"
   `include "rx_9600_5_no_2.sv"
   `include "rx_9600_6_no_2.sv"
   `include "rx_9600_7_no_2.sv"
   `include "rx_9600_8_no_2.sv"
   `include "rx_9600_5_even_2.sv"
   `include "rx_9600_6_even_2.sv"
   `include "rx_9600_7_even_2.sv"
   `include "rx_9600_8_even_2.sv"
   `include "rx_9600_5_odd_2.sv"
   `include "rx_9600_6_odd_2.sv"
   `include "rx_9600_7_odd_2.sv"
   `include "rx_9600_8_odd_2.sv"
   `include "rx_19200_5_no_1.sv"
   `include "rx_19200_6_no_1.sv"
   `include "rx_19200_7_no_1.sv"
   `include "rx_19200_8_no_1.sv"
   `include "rx_19200_5_even_1.sv"
   `include "rx_19200_6_even_1.sv"
   `include "rx_19200_7_even_1.sv"
   `include "rx_19200_8_even_1.sv"
   `include "rx_19200_5_odd_1.sv"
   `include "rx_19200_6_odd_1.sv"
   `include "rx_19200_7_odd_1.sv"
   `include "rx_19200_8_odd_1.sv"
   `include "rx_19200_5_no_2.sv"
   `include "rx_19200_6_no_2.sv"
   `include "rx_19200_7_no_2.sv"
   `include "rx_19200_8_no_2.sv"
   `include "rx_19200_5_even_2.sv"
   `include "rx_19200_6_even_2.sv"
   `include "rx_19200_7_even_2.sv"
   `include "rx_19200_8_even_2.sv"
   `include "rx_19200_5_odd_2.sv"
   `include "rx_19200_6_odd_2.sv"
   `include "rx_19200_7_odd_2.sv"
   `include "rx_19200_8_odd_2.sv"
   `include "rx_38400_5_no_1.sv"
   `include "rx_38400_6_no_1.sv"
   `include "rx_38400_7_no_1.sv"
   `include "rx_38400_8_no_1.sv"
   `include "rx_38400_5_even_1.sv"
   `include "rx_38400_6_even_1.sv"
   `include "rx_38400_7_even_1.sv"
   `include "rx_38400_8_even_1.sv"
   `include "rx_38400_5_odd_1.sv"
   `include "rx_38400_6_odd_1.sv"
   `include "rx_38400_7_odd_1.sv"
   `include "rx_38400_8_odd_1.sv"
   `include "rx_38400_5_no_2.sv"
   `include "rx_38400_6_no_2.sv"
   `include "rx_38400_7_no_2.sv"
   `include "rx_38400_8_no_2.sv"
   `include "rx_38400_5_even_2.sv"
   `include "rx_38400_6_even_2.sv"
   `include "rx_38400_7_even_2.sv"
   `include "rx_38400_8_even_2.sv"
   `include "rx_38400_5_odd_2.sv"
   `include "rx_38400_6_odd_2.sv"
   `include "rx_38400_7_odd_2.sv"
   `include "rx_38400_8_odd_2.sv"
   `include "rx_76800_5_no_1.sv"
   `include "rx_76800_6_no_1.sv"
   `include "rx_76800_7_no_1.sv"
   `include "rx_76800_8_no_1.sv"
   `include "rx_76800_5_even_1.sv"
   `include "rx_76800_6_even_1.sv"
   `include "rx_76800_7_even_1.sv"
   `include "rx_76800_8_even_1.sv"
   `include "rx_76800_5_odd_1.sv"
   `include "rx_76800_6_odd_1.sv"
   `include "rx_76800_7_odd_1.sv"
   `include "rx_76800_8_odd_1.sv"
   `include "rx_76800_5_no_2.sv"
   `include "rx_76800_6_no_2.sv"
   `include "rx_76800_7_no_2.sv"
   `include "rx_76800_8_no_2.sv"
   `include "rx_76800_5_even_2.sv"
   `include "rx_76800_6_even_2.sv"
   `include "rx_76800_7_even_2.sv"
   `include "rx_76800_8_even_2.sv"
   `include "rx_76800_5_odd_2.sv"
   `include "rx_76800_6_odd_2.sv"
   `include "rx_76800_7_odd_2.sv"
   `include "rx_76800_8_odd_2.sv"
   `include "rx_115200_5_no_1.sv"
   `include "rx_115200_6_no_1.sv"
   `include "rx_115200_7_no_1.sv"
   `include "rx_115200_8_no_1.sv"
   `include "rx_115200_5_even_1.sv"
   `include "rx_115200_6_even_1.sv"
   `include "rx_115200_7_even_1.sv"
   `include "rx_115200_8_even_1.sv"
   `include "rx_115200_5_odd_1.sv"
   `include "rx_115200_6_odd_1.sv"
   `include "rx_115200_7_odd_1.sv"
   `include "rx_115200_8_odd_1.sv"
   `include "rx_115200_5_no_2.sv"
   `include "rx_115200_6_no_2.sv"
   `include "rx_115200_7_no_2.sv"
   `include "rx_115200_8_no_2.sv"
   `include "rx_115200_5_even_2.sv"
   `include "rx_115200_6_even_2.sv"
   `include "rx_115200_7_even_2.sv"
   `include "rx_115200_8_even_2.sv"
   `include "rx_115200_5_odd_2.sv"
   `include "rx_115200_6_odd_2.sv"
   `include "rx_115200_7_odd_2.sv"
   `include "rx_115200_8_odd_2.sv"
   `include "rx_230400_5_no_1.sv"
   `include "rx_230400_6_no_1.sv"
   `include "rx_230400_7_no_1.sv"
   `include "rx_230400_8_no_1.sv"
   `include "rx_230400_5_even_1.sv"
   `include "rx_230400_6_even_1.sv"
   `include "rx_230400_7_even_1.sv"
   `include "rx_230400_8_even_1.sv"
   `include "rx_230400_5_odd_1.sv"
   `include "rx_230400_6_odd_1.sv"
   `include "rx_230400_7_odd_1.sv"
   `include "rx_230400_8_odd_1.sv"
   `include "rx_230400_5_no_2.sv"
   `include "rx_230400_6_no_2.sv"
   `include "rx_230400_7_no_2.sv"
   `include "rx_230400_8_no_2.sv"
   `include "rx_230400_5_even_2.sv"
   `include "rx_230400_6_even_2.sv"
   `include "rx_230400_7_even_2.sv"
   `include "rx_230400_8_even_2.sv"
   `include "rx_230400_5_odd_2.sv"
   `include "rx_230400_6_odd_2.sv"
   `include "rx_230400_7_odd_2.sv"
   `include "rx_230400_8_odd_2.sv"


	 /*---------------------FULL-DUPLEX TEST----------------------*/
   `include "full_2400_5_no_1.sv"
   `include "full_2400_6_no_1.sv"
   `include "full_2400_7_no_1.sv"
   `include "full_2400_8_no_1.sv"
   `include "full_2400_5_even_1.sv"
   `include "full_2400_6_even_1.sv"
   `include "full_2400_7_even_1.sv"
   `include "full_2400_8_even_1.sv"
   `include "full_2400_5_odd_1.sv"
   `include "full_2400_6_odd_1.sv"
   `include "full_2400_7_odd_1.sv"
   `include "full_2400_8_odd_1.sv"
   `include "full_2400_5_no_2.sv"
   `include "full_2400_6_no_2.sv"
   `include "full_2400_7_no_2.sv"
   `include "full_2400_8_no_2.sv"
   `include "full_2400_5_even_2.sv"
   `include "full_2400_6_even_2.sv"
   `include "full_2400_7_even_2.sv"
   `include "full_2400_8_even_2.sv"
   `include "full_2400_5_odd_2.sv"
   `include "full_2400_6_odd_2.sv"
   `include "full_2400_7_odd_2.sv"
   `include "full_2400_8_odd_2.sv"
   `include "full_4800_5_no_1.sv"
   `include "full_4800_6_no_1.sv"
   `include "full_4800_7_no_1.sv"
   `include "full_4800_8_no_1.sv"
   `include "full_4800_5_even_1.sv"
   `include "full_4800_6_even_1.sv"
   `include "full_4800_7_even_1.sv"
   `include "full_4800_8_even_1.sv"
   `include "full_4800_5_odd_1.sv"
   `include "full_4800_6_odd_1.sv"
   `include "full_4800_7_odd_1.sv"
   `include "full_4800_8_odd_1.sv"
   `include "full_4800_5_no_2.sv"
   `include "full_4800_6_no_2.sv"
   `include "full_4800_7_no_2.sv"
   `include "full_4800_8_no_2.sv"
   `include "full_4800_5_even_2.sv"
   `include "full_4800_6_even_2.sv"
   `include "full_4800_7_even_2.sv"
   `include "full_4800_8_even_2.sv"
   `include "full_4800_5_odd_2.sv"
   `include "full_4800_6_odd_2.sv"
   `include "full_4800_7_odd_2.sv"
   `include "full_4800_8_odd_2.sv"
   `include "full_9600_5_no_1.sv"
   `include "full_9600_6_no_1.sv"
   `include "full_9600_7_no_1.sv"
   `include "full_9600_8_no_1.sv"
   `include "full_9600_5_even_1.sv"
   `include "full_9600_6_even_1.sv"
   `include "full_9600_7_even_1.sv"
   `include "full_9600_8_even_1.sv"
   `include "full_9600_5_odd_1.sv"
   `include "full_9600_6_odd_1.sv"
   `include "full_9600_7_odd_1.sv"
   `include "full_9600_8_odd_1.sv"
   `include "full_9600_5_no_2.sv"
   `include "full_9600_6_no_2.sv"
   `include "full_9600_7_no_2.sv"
   `include "full_9600_8_no_2.sv"
   `include "full_9600_5_even_2.sv"
   `include "full_9600_6_even_2.sv"
   `include "full_9600_7_even_2.sv"
   `include "full_9600_8_even_2.sv"
   `include "full_9600_5_odd_2.sv"
   `include "full_9600_6_odd_2.sv"
   `include "full_9600_7_odd_2.sv"
   `include "full_9600_8_odd_2.sv"
   `include "full_19200_5_no_1.sv"
   `include "full_19200_6_no_1.sv"
   `include "full_19200_7_no_1.sv"
   `include "full_19200_8_no_1.sv"
   `include "full_19200_5_even_1.sv"
   `include "full_19200_6_even_1.sv"
   `include "full_19200_7_even_1.sv"
   `include "full_19200_8_even_1.sv"
   `include "full_19200_5_odd_1.sv"
   `include "full_19200_6_odd_1.sv"
   `include "full_19200_7_odd_1.sv"
   `include "full_19200_8_odd_1.sv"
   `include "full_19200_5_no_2.sv"
   `include "full_19200_6_no_2.sv"
   `include "full_19200_7_no_2.sv"
   `include "full_19200_8_no_2.sv"
   `include "full_19200_5_even_2.sv"
   `include "full_19200_6_even_2.sv"
   `include "full_19200_7_even_2.sv"
   `include "full_19200_8_even_2.sv"
   `include "full_19200_5_odd_2.sv"
   `include "full_19200_6_odd_2.sv"
   `include "full_19200_7_odd_2.sv"
   `include "full_19200_8_odd_2.sv"
   `include "full_38400_5_no_1.sv"
   `include "full_38400_6_no_1.sv"
   `include "full_38400_7_no_1.sv"
   `include "full_38400_8_no_1.sv"
   `include "full_38400_5_even_1.sv"
   `include "full_38400_6_even_1.sv"
   `include "full_38400_7_even_1.sv"
   `include "full_38400_8_even_1.sv"
   `include "full_38400_5_odd_1.sv"
   `include "full_38400_6_odd_1.sv"
   `include "full_38400_7_odd_1.sv"
   `include "full_38400_8_odd_1.sv"
   `include "full_38400_5_no_2.sv"
   `include "full_38400_6_no_2.sv"
   `include "full_38400_7_no_2.sv"
   `include "full_38400_8_no_2.sv"
   `include "full_38400_5_even_2.sv"
   `include "full_38400_6_even_2.sv"
   `include "full_38400_7_even_2.sv"
   `include "full_38400_8_even_2.sv"
   `include "full_38400_5_odd_2.sv"
   `include "full_38400_6_odd_2.sv"
   `include "full_38400_7_odd_2.sv"
   `include "full_38400_8_odd_2.sv"
   `include "full_76800_5_no_1.sv"
   `include "full_76800_6_no_1.sv"
   `include "full_76800_7_no_1.sv"
   `include "full_76800_8_no_1.sv"
   `include "full_76800_5_even_1.sv"
   `include "full_76800_6_even_1.sv"
   `include "full_76800_7_even_1.sv"
   `include "full_76800_8_even_1.sv"
   `include "full_76800_5_odd_1.sv"
   `include "full_76800_6_odd_1.sv"
   `include "full_76800_7_odd_1.sv"
   `include "full_76800_8_odd_1.sv"
   `include "full_76800_5_no_2.sv"
   `include "full_76800_6_no_2.sv"
   `include "full_76800_7_no_2.sv"
   `include "full_76800_8_no_2.sv"
   `include "full_76800_5_even_2.sv"
   `include "full_76800_6_even_2.sv"
   `include "full_76800_7_even_2.sv"
   `include "full_76800_8_even_2.sv"
   `include "full_76800_5_odd_2.sv"
   `include "full_76800_6_odd_2.sv"
   `include "full_76800_7_odd_2.sv"
   `include "full_76800_8_odd_2.sv"
   `include "full_115200_5_no_1.sv"
   `include "full_115200_6_no_1.sv"
   `include "full_115200_7_no_1.sv"
   `include "full_115200_8_no_1.sv"
   `include "full_115200_5_even_1.sv"
   `include "full_115200_6_even_1.sv"
   `include "full_115200_7_even_1.sv"
   `include "full_115200_8_even_1.sv"
   `include "full_115200_5_odd_1.sv"
   `include "full_115200_6_odd_1.sv"
   `include "full_115200_7_odd_1.sv"
   `include "full_115200_8_odd_1.sv"
   `include "full_115200_5_no_2.sv"
   `include "full_115200_6_no_2.sv"
   `include "full_115200_7_no_2.sv"
   `include "full_115200_8_no_2.sv"
   `include "full_115200_5_even_2.sv"
   `include "full_115200_6_even_2.sv"
   `include "full_115200_7_even_2.sv"
   `include "full_115200_8_even_2.sv"
   `include "full_115200_5_odd_2.sv"
   `include "full_115200_6_odd_2.sv"
   `include "full_115200_7_odd_2.sv"
   `include "full_115200_8_odd_2.sv"
   `include "full_230400_5_no_1.sv"
   `include "full_230400_6_no_1.sv"
   `include "full_230400_7_no_1.sv"
   `include "full_230400_8_no_1.sv"
   `include "full_230400_5_even_1.sv"
   `include "full_230400_6_even_1.sv"
   `include "full_230400_7_even_1.sv"
   `include "full_230400_8_even_1.sv"
   `include "full_230400_5_odd_1.sv"
   `include "full_230400_6_odd_1.sv"
   `include "full_230400_7_odd_1.sv"
   `include "full_230400_8_odd_1.sv"
   `include "full_230400_5_no_2.sv"
   `include "full_230400_6_no_2.sv"
   `include "full_230400_7_no_2.sv"
   `include "full_230400_8_no_2.sv"
   `include "full_230400_5_even_2.sv"
   `include "full_230400_6_even_2.sv"
   `include "full_230400_7_even_2.sv"
   `include "full_230400_8_even_2.sv"
   `include "full_230400_5_odd_2.sv"
   `include "full_230400_6_odd_2.sv"
   `include "full_230400_7_odd_2.sv"
   `include "full_230400_8_odd_2.sv"

	/*-----------INTERRUPT-------------*/
	`include "parity_error_en.sv"
	`include "parity_error_dis.sv"
	`include "tx_fifo_empty_en.sv"
	`include "tx_fifo_empty_dis.sv"
	`include "tx_fifo_full_en.sv"
	`include "tx_fifo_full_dis.sv"
	`include "rx_fifo_empty_en.sv"
	`include "rx_fifo_empty_dis.sv"
	`include "rx_fifo_full_en.sv"
	`include "rx_fifo_full_dis.sv"

	/*-----------ERROR INJECTION TEST-------------*/
	`include "data_bits_mismatch.sv"
	`include "baudrate_mismatch.sv"
	`include "parity_mismatch.sv"
	`include "stop_bits_mismatch.sv"
	
	/*-----------ERROR HANDLING-------------*/
	`include "write_tx_fifo_full.sv"
	`include "access_rsvd.sv"	


	/*-----------DYNAMIC RECONFIG - TX-------------*/
	`include "tx_baudrate_reconfig.sv"
	`include "tx_data_bits_reconfig.sv"
	`include "tx_parity_reconfig.sv"
	`include "tx_stop_bits_reconfig.sv"

	/*-----------DYNAMIC RECONFIG - RX-------------*/
	`include "rx_baudrate_reconfig.sv"
	`include "rx_data_bits_reconfig.sv"
	`include "rx_parity_reconfig.sv"
	`include "rx_stop_bits_reconfig.sv"

	/*-----------DYNAMIC RECONFIG - FULL-------------*/
	`include "full_baudrate_reconfig.sv"
	`include "full_data_bits_reconfig.sv"
	`include "full_parity_reconfig.sv"
	`include "full_stop_bits_reconfig.sv" 
endpackage
